-- This file is automatically generate and will be overwriten the next time the script runs




library ieee;
use ieee.std_logic_1164.all;

package RAM_DATA is

constant RAM0 : string := "00010111,00010011,11101111,01100011,10110111,10000011,00010011,00100011,00100011,"&
"00110111,00100011,00100011,10110111,00100011,00100011,00100011,00100011,10010011,"&
"00100011,10010011,00100011,00110111,10010011,00010011,10000011,01100011,10000011,"&
"00000011,10000011,00000011,10000011,00000011,10000011,00010011,01100111,10000011,"&
"00100011,00000011,10000011,01100011,10000011,00000011,10000011,10110011,10110011,"&
"10110011,00100011,10000011,00100011,10000011,11100011,00000011,00000011,10010011,"&
"11101111,00110011,00100011,00000011,10010011,11101111,00100011,01101111,10000011,"&
"00000011,10000011,10110011,01101111,00110111,10000011,10010011,11100011,10110111,"&
"00100011,01100111,01100011,00000011,00100011,00000011,00010011,00100011,01100111,"&
"01100011,00010011,01101111,01100111,00010011,00100011,10110111,10010011,00100011,"&
"00100011,00100011,00100011,00100011,00100011,00100011,00100011,00100011,00100011,"&
"10010011,00010011,10010011,00100011,10000011,01100011,00010011,10010011,11101111,"&
"10000011,00000011,10000011,00000011,10000011,00000011,10000011,00000011,10000011,"&
"00000011,10000011,00010011,00010011,01100111,10010011,01100011,00010011,11101111,"&
"00010011,01101111,00000011,10010011,01100011,00010011,00010011,10000011,10010011,"&
"00010011,10010011,10010011,01100011,00010011,10010011,01101111,00010011,01101111,"&
"10010011,00110011,00010011,00110011,00010011,00010011,10000011,00010011,10010011,"&
"10010011,11100011,10000011,10010011,01100011,00010011,10000011,10010011,01100011,"&
"01100011,10010011,01100011,10010011,11100011,10000011,00010011,00010011,11101111,"&
"10010011,01101111,10010011,01100011,10010011,01100011,10010011,11100011,10000011,"&
"00010011,01100011,10110111,10010011,10000011,01100011,01100011,01100011,10010011,"&
"01101111,00010011,11101111,10010011,00010011,01101111,10010011,00010011,11101111,"&
"00010011,01101111,00000011,00010011,10010011,01100011,10010011,00100011,10010011,"&
"00110011,01100011,00010011,10010011,11100011,10010011,10110011,10000011,00010011,"&
"11101111,01101111,00000011,10010011,00010011,01101111,00000011,10010011,10010011,"&
"11100011,10010011,00010011,00110011,11101111,00010011,00010011,10010011,10010011,"&
"10010011,00010011,11101111,10000011,10010011,10010011,00110011,10000011,00010011,"&
"10010011,00100011,11101111,10010011,00010011,11100011,01101111,10010011,00010011,"&
"11101111,00010011,01101111,10110111,00000011,00010011,01100111,00110111,10000011,"&
"10010011,11100011,10110111,00000011,01100111,10010011,01100011,01100111,00110011,"&
"10000011,00110011,10010011,00100011,01101111,00110011,10010011,01100011,01100111,"&
"10010011,10100011,01101111,00010011,00100011,00100011,00100011,00100011,00100011,"&
"00100011,00100011,00100011,00100011,00000011,10010011,00010011,00010011,10010011,"&
"01100011,00010011,10010011,00000011,10010011,01100011,00000011,10010011,01100011,"&
"00010011,00010011,00010011,00010011,10010011,10010011,00010011,10000011,10010011,"&
"01100011,00010011,10010011,01100011,00010011,01100011,10010011,10010011,00010011,"&
"00100011,11101111,00110011,00000011,01100011,01100011,00100011,01100011,00110011,"&
"10000011,00000011,10000011,00000011,10000011,00000011,10000011,00000011,10000011,"&
"00010011,01100111,00010011,01101111,00010011,00100011,00100011,00100011,00100011,"&
"00100011,00010011,00010011,10010011,10010011,11101111,01100011,01100011,01100011,"&
"00010011,01101111,01100011,00100011,00010011,10000011,00000011,10000011,00000011,"&
"10000011,00010011,01100111,10010011,10100011,01101111,00010011,00100011,00100011,"&
"10010011,00010011,00010011,00100011,00100011,00100011,00100011,00100011,00100011,"&
"00100011,11101111,10000011,00010011,01100111,00010011,00100011,00100011,00100011,"&
"00100011,00100011,00100011,00100011,00100011,00100011,00100011,00100011,00010011,"&
"00010011,00010011,10110111,00110111,10010011,10010011,00110111,10010011,10110011,"&
"01100011,10000011,00000011,10000011,00000011,10000011,00000011,10000011,00000011,"&
"10000011,00000011,10000011,00010011,00010011,01100111,10010011,00010011,11101111,"&
"10010011,10110011,10000011,00010011,11101111,01100011,00010011,11101111,10010011,"&
"11100011,00010011,11101111,10010011,10110011,00000011,10010011,10010011,01100011,"&
"10010011,11101111,11100011,00010011,11101111,00010011,01101111,00010011,01101111,"&
"10010011,01100011,00010011,01100111,00010011,01100011,10110011,00010011,10010011,"&
"01101111,10010011,00010011,01100011,10010011,01100011,01100011,10010011,01100011,"&
"01100011,10010011,00010011,01100111,10010011,00010011,01101111,01100011,00110011,"&
"10110011,00010011,10010011,01101111,00010011,01101111,00010011,01101111,10110111,"&
"00010011,00100011,00100011,10110111,00000011,00010011,00100011,00000011,00010011,"&
"00100011,00110111,10000011,10010011,00100011,01100111,10110111,00000011,10110111,"&
"10010011,01100011,00110111,00010011,00010011,10110111,00110111,00100011,11101111,"&
"10000011,00010011,00110111,00010011,01100111,01100111,10110111,00110111,00010011,"&
"10010011,00010011,00100011,00100011,00100011,00100011,00100011,00100011,00100011,"&
"00100011,00100011,00100011,00100011,10110111,11101111,00110111,00010011,00110111,"&
"10110111,00110111,10110111,00010011,11101111,10110111,00010011,11101111,10110111,"&
"00010011,11101111,00010011,11101111,00010011,11101111,00010011,11101111,00110111,"&
"00010011,11101111,00110111,00010011,11101111,11101111,10010011,11101111,10010011,"&
"01100011,01100011,10010011,01100011,01100011,10010011,01100011,10010011,11100011,"&
"01100011,00110111,00010011,11101111,01101111,10010011,01100011,10010011,11100011,"&
"00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,11101111,"&
"10010011,00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,"&
"11101111,10010011,00010011,11101111,01101111,10010011,01100011,01100011,10010011,"&
"01100011,10010011,11100011,00110111,00010011,11101111,00010011,11101111,10010011,"&
"00010011,00010011,11101111,10000011,00110111,00010011,11101111,01101111,10010011,"&
"01100011,10010011,11100011,00110111,00010011,11101111,00010011,11101111,00010011,"&
"10010011,00010011,11101111,10010011,00110111,00010011,11101111,00010011,11101111,"&
"00010011,10010011,00010011,11101111,00100011,01101111,00110111,00010011,11101111,"&
"10110111,00110111,01101111,00110111,00010011,11101111,10110111,00110111,01101111,"&
"00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,11101111,"&
"10010011,00010011,00110111,10010011,00010011,11101111,11101111,00010011,00010011,"&
"10110111,10110011,00100011,00010011,11101111,01100011,11101111,10010011,00010011,"&
"01100011,00010011,11101111,00010011,01101111,00010011,11100011,00010011,01101111,"&
"00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,11101111,"&
"00010011,00110111,00010011,11101111,00010011,11100111,01101111,00110111,00010011,"&
"11101111,11101111,00010011,10010011,11100011,10010011,10010011,00110111,10110111,"&
"00010011,00100011,10110011,10000011,00110011,00010011,00100011,11101111,00010011,"&
"01100011,00010011,11101111,10010011,11100011,00110111,10010011,00010011,01101111,"&
"00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,11101111,"&
"10010011,00110111,00010011,11101111,00010011,11101111,00010011,10010011,00010011,"&
"11101111,00010011,00110111,00010011,11101111,00010011,11101111,00010011,10010011,"&
"00010011,11101111,10010011,00010011,00010011,11101111,01101111,00010011,00100011,"&
"11101111,11101111,11101111,00001010,01111000,00100101,00100000,00100000,00111100,"&
"01001100,00110000,00110100,00111000,01100011,00000000,01010011,00100000,00110000,"&
"01001000,01001001,01010011,01100010,01101100,01100101,00100000,00000000,00001010,"&
"00100000,01110011,01100011,01010000,00100000,00100000,01001101,00001010,00100000,"&
"01110101,01100001,01101001,01111001,00001010,00100000,01100010,00000000,00001010,"&
"00100000,01110000,01110010,01100101,01000101,01001111,00001010,00100000,01101000,"&
"01110101,00001010,00100000,01100110,00000000,00001010,00100000,01110010,00100000,"&
"01100100,00001010,00100000,01110111,01100101,01110010,00001010,00100000,01100101,"&
"01100100,00001010,01001101,01101100,01100101,00001010,01110010,00100000,01111000,"&
"00001010,01110100,00100000,00100000,01100001,01100001,01111000,01111000,00001010,"&
"00001010,01110100,00001010,01100100,00000000,00001010,01110100,01101111,01010000,"&
"00111111,00101101,00100101,01111001,00000000,00001010,01100111,00101000,00101001,"&
"00001010,01100101,01100101,00000000,00100101,00001010,00001010,01100100,01100101,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,";


constant RAM1 : string := "00000001,00000001,00000000,00000000,01000111,10100111,00000001,00100100,00100010,"&
"01100100,00100010,00100110,10000100,00101110,00101100,00101010,00100110,00001010,"&
"00100000,00001001,00100100,01001010,10000100,00000100,00100111,11100100,00100000,"&
"00100100,00100100,00101001,00101001,00101010,00101010,00000001,10000000,00100111,"&
"00100000,00100111,00100111,01111110,00100111,00100111,00100110,10000111,10000111,"&
"10000111,00100100,00100111,00100010,00100111,11111100,00100101,00101001,00000101,"&
"00000000,00000101,00100110,00100101,00000101,00000000,00100100,11110000,00100111,"&
"00100111,00100110,10000111,11110000,00000111,00100111,11110111,10011100,01000111,"&
"10100000,10000000,00001110,00100111,00000000,00100111,00000111,00100000,10000000,"&
"10000110,10000101,11110000,10000000,00000001,00101010,00011010,10000111,00101110,"&
"00101000,00100110,00100110,00100100,00100010,00100000,00101100,00100100,00100010,"&
"00001001,10001011,00001011,00100110,01000101,10010100,10000101,00000101,11110000,"&
"00100000,00100100,00100100,00101001,00101001,00101010,00101010,00101011,00101011,"&
"00101100,00101100,00000101,00000001,10000000,00000111,10001010,10000101,11110000,"&
"00001011,11110000,01001010,00000111,00001000,00001011,00001010,01000111,00000110,"&
"00000100,10000111,11110111,11100010,00000100,00000101,00000000,00001011,11110000,"&
"00010111,10000100,00010100,00000100,00000100,00001011,01000110,00000101,10000111,"&
"11110111,11111100,01000110,00000111,10010100,00001011,01000111,00000110,10001010,"&
"11100110,00000110,10001000,00000110,10010000,11000101,10000100,10000101,11110000,"&
"00001011,11110000,00000110,10001000,00000110,10000000,00000110,10011000,10100100,"&
"10001001,10010110,00010111,10000100,11000101,10000100,00011000,01000000,00001011,"&
"11110000,10000101,11110000,10000100,00000100,11110000,00000101,10000101,11110000,"&
"00000100,11110000,10101001,00001100,10001011,00011010,00000111,00001000,00000100,"&
"00000100,01000100,00000100,10000100,10000110,00000111,10000111,11000101,10000101,"&
"11110000,11110000,10101001,10001011,00001100,11110000,10101001,10000100,10001011,"&
"01010110,00000101,10000101,00001001,11110000,00000100,00001100,00001100,00000100,"&
"00000101,00000101,00000000,00100111,00000101,00001010,10000101,01000110,00000101,"&
"10000100,10000000,00000000,10001100,00001001,11110100,11110000,00000101,10000101,"&
"11110000,00000100,11110000,00000111,10100101,01110101,10000000,00000111,00100111,"&
"11110111,10001100,01000111,10100101,10000000,00000111,00010100,10000000,10000111,"&
"01000110,00000111,10000111,00000000,11110000,00000110,00000111,10010100,10000000,"&
"10000111,10001111,11110000,00000001,00101100,00100110,00100100,00101110,00101010,"&
"00101000,00100010,00100000,00101110,01000111,00000111,00000100,10001010,00001001,"&
"00010110,00000100,00001001,01000111,00000111,00011100,01000111,00000111,00010110,"&
"00000100,00000110,00001011,00000101,00001011,00001010,00001001,01000111,10000100,"&
"11111110,10000111,10000100,11111000,10000111,11100010,10000100,00000101,00000101,"&
"00100110,00000000,00000101,00100110,00010000,00000100,00100000,10000100,00000101,"&
"00100000,00100100,00100100,00101001,00101001,00101010,00101010,00101011,00101011,"&
"00000001,10000000,00000100,11110000,00000001,00101100,00101010,00101000,00100110,"&
"00101110,00000100,00001001,00000100,00001001,11110000,00001100,01011000,10011000,"&
"00000101,00000000,10010100,10000000,00000101,00100000,00100100,00100100,00101001,"&
"00101001,00000001,10000000,10000100,10001111,11110000,00000001,00100010,00100100,"&
"00000101,00000110,00000101,00101110,00100110,00101000,00101010,00101100,00101110,"&
"00100110,11110000,00100000,00000001,10000000,00000001,00100100,00100000,00101110,"&
"00101100,00101010,00101000,00100110,00100100,00100010,00100110,00100010,00001001,"&
"10001010,00000100,00011010,00011011,00001011,00001001,00011100,00001100,00000111,"&
"11101110,00100000,00100100,00100100,00101001,00101001,00101010,00101010,00101011,"&
"00101011,00101100,00101100,00000101,00000001,10000000,00000101,10000101,11110000,"&
"00000100,00000111,11000101,00000101,11110000,10010110,00000101,11110000,10000100,"&
"10010000,00000101,11110000,00000100,00000111,11000101,00000111,11110111,11100000,"&
"10000100,11110000,10010010,00000101,11110000,00000100,11110000,00000101,11110000,"&
"00000111,10010110,10000101,10000000,11110111,00000100,10000111,00010101,11010101,"&
"11110000,00000111,00000111,11111000,10000111,10001000,11011110,00000111,00010000,"&
"00000100,00000111,10000101,10000000,10010101,00010111,11110000,01100110,00000101,"&
"11100111,01010111,11010101,11110000,00000110,11110000,00000110,11110000,01000111,"&
"00000111,10101000,10100000,01000111,10100111,01100111,10100000,10100111,01110111,"&
"10100000,01000111,00100111,11100111,00100000,10000000,00000111,10100111,01110111,"&
"10000111,00011010,00100110,00000001,00000110,00000101,00000101,00100110,11110000,"&
"00100000,00000101,00000011,00000001,00000000,10000000,00010101,00010101,00000001,"&
"10000101,00000101,00101100,00101010,00101000,00100100,00100010,00100000,00101110,"&
"00100110,00101110,00101100,00101010,00000100,11110000,00001001,00000100,00011010,"&
"00011010,00011011,00010111,10000101,11110000,00010111,10000101,11110000,00010111,"&
"10000101,11110000,00000101,11110000,10000101,11110000,00000101,11110000,00010101,"&
"00000101,11110000,00010101,00000101,11110000,11110000,00001011,11110000,00000111,"&
"10001010,11000000,00000111,10000000,11000100,00000111,10000010,00000111,10011110,"&
"00011100,00010101,00000101,11110000,11110000,00000111,10000100,00000111,10011100,"&
"00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,11110000,"&
"00001011,00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,"&
"11110000,00000101,10000101,11110000,11110000,00000111,10001010,11000110,00000111,"&
"10001110,00000111,10010000,00010101,00000101,11110000,00000101,11110000,00000101,"&
"00000110,00000101,11110000,01000101,00010101,00000101,11110000,11110000,00000111,"&
"10001110,00000111,10011100,00010101,00000101,11110000,00000101,11110000,00000110,"&
"00000101,00000101,11110000,00001011,00010101,00000101,11110000,00000101,11110000,"&
"00000110,00000101,00000101,11110000,10000000,11110000,00010101,00000101,11110000,"&
"00000100,00001001,11110000,00010101,00000101,11110000,00000100,00001001,11110000,"&
"00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,11110000,"&
"00000100,00001001,00010101,10000101,00000101,11110000,11110000,00001100,00000100,"&
"11011011,10000111,10000000,10001100,11110000,00000010,11110000,01110111,00001100,"&
"10010110,00000101,11110000,00000100,11110000,00001100,00011010,00000100,00000000,"&
"00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,11110000,"&
"00001001,00010101,00000101,11110000,00000101,00000000,11110000,00010101,00000101,"&
"11110000,11110000,01110101,00000111,00010100,01011011,00001001,00001100,00001100,"&
"10010111,00000000,10000110,10100110,00000111,00000101,00100000,11110000,11110111,"&
"00010110,00000101,11110000,10001001,11010110,00010101,00000101,00000101,11110000,"&
"00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,11110000,"&
"00001011,00010101,00000101,11110000,00000101,11110000,00000110,00000101,00000101,"&
"11110000,00001100,00010101,00000101,11110000,00000101,11110000,00000110,00000101,"&
"00000101,11110000,01110101,00000110,10000101,11110000,11110000,00000001,00100110,"&
"11110000,11110000,11110000,00100101,00100000,00110000,00000000,01111100,01001110,"&
"00111110,00110001,00110101,00111001,01100100,00000000,01100101,00110001,00110001,"&
"01000110,01010011,01101111,01101111,01101111,01110010,00100101,00000000,01011011,"&
"01100101,01100101,01110100,01001101,01100101,01010011,00000000,01011011,01010101,"&
"01110000,01100100,01101110,00000000,01011011,01000010,01101111,00000000,01011011,"&
"00100000,01110010,01100001,01111000,01000101,01001101,01011011,00100000,01100101,"&
"01101101,01011011,00100000,01101001,00000000,01011011,00100000,01100101,01110111,"&
"00000000,01011011,00100000,01110010,00100000,01100100,01010011,01110011,01100011,"&
"00000000,01010011,00100000,01100101,01100100,01100001,01100101,00101000,00101001,"&
"01110111,01101001,01100110,01100010,01110010,01110100,00100101,00101110,00000000,"&
"01100010,00001010,01101110,01100001,00000000,01110111,01100101,00100000,01010010,"&
"00001010,00101101,01100100,01110100,00000000,01101100,01110100,01101000,00111010,"&
"01100010,00100000,01111000,00000000,00110000,00000000,01110111,00100000,01111000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,";


constant RAM2 : string := "00000000,11000001,00010000,00000000,00000010,00000111,00000001,10000001,11110001,"&
"00000000,10010001,00000001,01111101,00110001,01000001,01010001,00010001,01110100,"&
"00100001,00000101,00000001,00000010,00000100,10000100,11000001,00110111,11000001,"&
"10000001,01000001,00000001,11000001,10000001,01000001,00000001,00000000,00001010,"&
"11110001,00000001,01000001,11110111,00000001,01000001,10000001,11010111,10010111,"&
"11100111,11110001,00000001,11110001,10000001,11111010,10000001,11000001,00000100,"&
"00000000,00100101,10100001,10000001,00000100,01000000,10100001,11011111,00000001,"&
"01000001,10000001,11010111,11011111,00000011,00000111,00100111,00000111,00000011,"&
"10100111,00000000,00000101,00000101,10110111,00000101,00010111,11100101,00000000,"&
"00000101,00000101,00011111,00000000,00000001,01010001,00000000,10001010,00110001,"&
"01100001,01110001,00010001,10000001,10010001,00100001,01000001,10000001,10010001,"&
"00000101,00000101,00000110,11110001,00001011,00000101,00001001,00000000,11011111,"&
"11000001,10000001,01000001,00000001,11000001,10000001,01000001,00000001,11000001,"&
"10000001,01000001,00000000,00000001,00000000,01010000,11110101,00001001,01011111,"&
"00011011,00011111,00011011,00000000,11111010,00011011,00000000,00001011,10010000,"&
"11110000,00000111,11110111,11110110,00000000,10010000,01000000,00101011,10011111,"&
"00100100,10000111,00010100,11010100,00000100,00000101,00001011,00011011,00000110,"&
"11110111,11110101,00001011,11000000,11110110,00011011,00001011,01000000,11010111,"&
"11110110,10000000,11010111,00110000,11010111,00001011,01001011,00001001,00011111,"&
"00000100,10011111,01010000,11010111,10000000,11010111,00110000,11010111,00001011,"&
"01001011,00000100,00000000,00000111,00000100,00000101,00000100,10000000,00001001,"&
"01011111,00001001,11011111,00010100,11110100,10011111,00001010,00001001,01011111,"&
"11110100,00011111,00001011,00000000,01001011,00001001,00000000,11110001,00010000,"&
"10010100,10000000,11110000,11110100,10000100,00000001,10010111,00000111,00001001,"&
"10011111,01011111,00001011,01001011,10100000,10011111,00001011,01001011,00000100,"&
"00001001,11010000,00001001,00100000,01011111,11110100,10100000,00000001,00000000,"&
"00001100,00001001,00000000,11000001,00001100,00001001,10100111,00000101,00001001,"&
"00010100,11011100,01000000,00011100,00000101,10001010,10011111,00001010,00001001,"&
"10011111,11110100,10011111,00000011,00000111,00010101,00000000,00000011,00000111,"&
"00010111,00000111,00000011,00000111,00000000,00000000,11110110,00000000,11110101,"&
"00000111,11110101,00010111,11010111,01011111,11000101,00000101,11000111,00000000,"&
"00010111,10110111,00011111,00000001,10000001,00110001,01000001,00010001,10010001,"&
"00100001,01010001,01100001,01110001,00000101,11010000,00000101,00000101,00000000,"&
"11110111,00010101,00010000,00000100,00000000,11110111,00010100,10000000,11110111,"&
"00100100,00000000,10010100,00000000,10010000,10010000,00010100,11111001,00000111,"&
"10011011,11110111,10010111,11101010,11110111,11101010,10010111,00000101,00000110,"&
"11000001,10000000,10010101,11000001,00101011,00001010,10001010,00001001,10100000,"&
"11000001,10000001,01000001,00000001,11000001,10000001,01000001,00000001,11000001,"&
"00000001,00000000,00001001,11011111,00000001,10000001,10010001,00100001,00110001,"&
"00010001,00000101,11110101,00000101,10100000,11011111,00110101,00000101,10000100,"&
"00000000,00000000,00100100,00000100,00000100,11000001,10000001,01000001,00000001,"&
"11000001,00000001,00000000,00010100,10100100,10011111,00000001,10110001,11000001,"&
"00000101,01000001,00000000,00010001,11010001,11100001,11110001,00000001,00010001,"&
"11000001,01011111,11000001,00000001,00000000,00000001,10000001,00100001,00110001,"&
"01000001,01010001,01100001,01110001,10000001,10010001,00010001,10010001,00000101,"&
"00000101,00000101,00000000,00000000,01110000,00000000,00000000,11100000,00100100,"&
"01000111,11000001,10000001,01000001,00000001,11000001,10000001,01000001,00000001,"&
"11000001,10000001,01000001,00000000,00000001,00000000,00000100,11001010,00011111,"&
"00000000,10010100,00000111,01001011,11011111,01110100,00000000,00011111,00010100,"&
"00110100,11001100,00011111,00000000,10010100,00000111,00000101,11110111,11111100,"&
"00010100,00011111,00110100,11000000,01011111,00000100,01011111,11100000,00011111,"&
"00000000,00000101,00000111,00000000,00010101,00000111,10100111,00010101,00010101,"&
"00011111,00010000,00010000,10100101,11110111,00000111,00000101,00000000,00000111,"&
"00000110,00000101,00000111,00000000,00010101,00010111,00011111,10110101,10110101,"&
"11100111,00010111,00010101,11011111,00000000,10011111,00010000,00011111,00000011,"&
"00100000,11100111,00000111,00000001,00000111,01000111,11100111,00000111,01110111,"&
"11100111,00000000,00000111,00000111,11110111,00000000,00000000,00000111,00000000,"&
"00010111,11110111,00000000,00000001,00000110,00000000,00000000,00010001,01011111,"&
"11000001,00000000,00000000,00000001,00000011,00000000,00000000,00000000,00000001,"&
"11000101,10000101,10000001,10010001,00100001,01000001,01010001,01100001,00010001,"&
"00110001,01110001,10000001,10010001,00000000,10011111,00000000,00000000,00000000,"&
"00000000,00000000,00000000,10000111,10011111,00000000,10000111,11011111,00000000,"&
"00000111,00011111,00001010,10011111,11001010,00011111,11001011,10011111,00000000,"&
"11000101,11011111,00000000,00000101,00011111,11011111,00000101,01011111,01010000,"&
"11111011,01110111,01010000,11111011,01110111,00100000,11111011,00000000,11111011,"&
"00000100,00000000,00000101,11011111,10011111,00100000,11111011,01000000,11111011,"&
"00000000,01000101,11011111,00000001,00011111,00000000,00000000,00000001,00011111,"&
"00000101,00000000,00000101,01011111,00000001,10011111,00000000,00000000,00000001,"&
"10011111,00000101,00001011,01011111,11011111,00110000,11111011,01110111,01100000,"&
"11111011,00100000,11111011,00000000,01000101,01011111,00000001,10011111,00000000,"&
"00000000,00000001,10011111,00000101,00000000,00000101,11011111,10011111,01010000,"&
"11111011,01110000,11111011,00000000,01000101,11011111,00000001,00011111,00000000,"&
"00000000,00000001,00011111,00000101,00000000,10000101,01011111,00000001,10011111,"&
"00000000,00000000,00000001,10011111,10101011,01011111,00000000,01000101,10011111,"&
"00000000,00000000,11011111,00000000,01000101,00011111,00000000,00000000,01011111,"&
"00000000,01000101,10011111,00000001,11011111,00000000,00000000,00000001,11011111,"&
"00000101,00000101,00000000,00000100,01000101,10011111,01011111,00000101,00000000,"&
"00000011,10000100,10000111,00001011,10011111,00000101,00011111,11110100,00000101,"&
"00000111,00110000,11001111,00010100,00011111,11111100,00001100,00010100,10000000,"&
"00000000,01000101,10011111,00000001,11011111,00000000,00000000,00000001,11011111,"&
"00000101,00000000,10000101,00011111,00000000,00001001,01011111,00000000,11000101,"&
"10011111,01011111,11110101,10010000,11110101,00100100,00000000,10000000,00000000,"&
"00101001,00001100,11100100,00000110,10010111,01010000,11010111,11001111,11111001,"&
"00000111,00110000,10001111,00011001,00111011,00000000,00000100,00000101,01011111,"&
"00000000,01000101,01011111,00000001,10011111,00000000,00000000,00000001,10011111,"&
"00000101,00000000,00000101,11011111,00000001,00011111,00000000,00000000,00000001,"&
"00011111,00000101,00000000,00000101,01011111,00000001,10011111,00000000,00000000,"&
"00000001,10011111,11110101,00001100,00001011,11001111,10011111,00000001,00010001,"&
"10011111,01011111,10011111,00110000,00000000,00110010,00000000,00000000,01010101,"&
"00000000,00110010,00110110,01100001,01100101,00000000,01110000,00100000,00111001,"&
"00101101,01000011,01000011,01101111,01100001,00100000,01110011,00000000,01110011,"&
"01011101,01101100,00100000,00100000,01111000,01010010,00000000,01110101,01011101,"&
"01101100,00100000,01100001,00000000,01100010,01011101,01101111,00000000,01010000,"&
"01011101,01101111,01101101,01110100,01010000,00000000,01100100,01011101,01111000,"&
"01110000,01100110,01011101,01101100,00000000,01110010,01011101,01100001,01101111,"&
"00000000,01110111,01011101,01101001,01110111,00001010,01010000,01100101,01110100,"&
"00000000,01010010,01110011,01100011,00000000,01100100,01110011,01101000,00111010,"&
"01100001,01101110,01101111,01101001,01111001,00100000,00110000,00101110,00000000,"&
"01101111,00000000,01101111,01110100,00000000,01110010,00100000,01000101,01001111,"&
"00000000,00111110,00100000,01100101,00000000,01100101,01101000,01100101,00000000,"&
"01111001,00101000,00101001,00000000,00111000,00000000,01101111,00101000,00101001,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,";


constant RAM3 : string := "01010000,11111111,01000101,00000000,11100001,00000000,11111101,00000010,00000000,"&
"00000000,00000010,00000000,00000001,00000001,00000001,00000001,00000010,00011010,"&
"00000011,00000000,00000000,11100001,10000100,00011010,00000000,00000011,00000010,"&
"00000010,00000010,00000010,00000001,00000001,00000001,00000011,00000000,00000000,"&
"00000000,00000000,00000000,00000100,00000000,00000000,00000000,00000000,00000000,"&
"01000000,00000000,00000000,00000000,00000000,11111000,00000000,00000000,00000000,"&
"01101101,00000001,00000000,00000000,00000000,01101100,00000000,11110110,00000000,"&
"00000000,00000000,00000000,11111010,11100001,01000000,00000000,11111110,11100001,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,11111100,00000000,11111011,00000011,00000000,11001000,00000011,"&
"00000011,00000011,00000100,00000100,00000100,00000101,00000011,00000011,00000011,"&
"00000000,00000000,00000000,00000000,00000000,00000100,00000000,00000000,11110111,"&
"00000100,00000100,00000100,00000100,00000011,00000011,00000011,00000011,00000010,"&
"00000010,00000010,00000000,00000101,00000000,00000010,00000000,00000000,11110011,"&
"00000000,11111010,00000000,00000011,00000010,00000000,00000010,00000000,00000000,"&
"11111111,11111101,00001111,00000100,00000000,00000000,00000010,00000000,11111101,"&
"00000000,00000000,00000000,00000000,11111101,00000000,00000000,00000000,11111101,"&
"00001111,11111100,00000000,00000110,00000000,00000000,00000000,00000110,00001110,"&
"00000010,00000101,00001000,00000110,11110110,00000000,00000000,00000000,11101000,"&
"00000000,11110100,00000111,00001010,00000111,00000110,00000111,11110010,00000000,"&
"00000000,00000000,00000000,11001000,00000000,00000000,00000000,00000010,00000000,"&
"11110000,00000000,11100010,00000000,11111111,11111101,00000000,00000000,11100001,"&
"11111111,11111101,00000000,00000001,00000000,00000110,00000011,00000000,00000000,"&
"01000000,00001010,11111111,11111111,11101010,00000001,00000000,00000000,00000000,"&
"11011100,11111110,00000000,00000000,00000000,11111011,00000000,00000000,00000000,"&
"11111110,00000010,00000000,01000001,11011001,11111111,00000000,00000001,00000000,"&
"00000000,00000000,01000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00111101,00000000,00000000,11111101,11110101,00000000,00000000,"&
"11010011,11111111,11110100,11100001,01000000,00000000,00000000,11100001,01000000,"&
"00000000,11111110,11100001,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,11111110,00000000,00000000,00000000,00000000,"&
"00000000,11111110,11111111,11111100,00000010,00000011,00000011,00000010,00000010,"&
"00000011,00000011,00000011,00000001,00000000,00000010,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000011,00000000,00000000,00000111,00000000,"&
"00000000,00000001,00000000,00000000,00000000,00000001,00000000,11111111,11111101,"&
"00000000,11111011,11111100,00000000,11111001,00000010,11111010,00000000,00000000,"&
"00000000,00100001,00000000,00000000,00000101,00000000,00000000,00000000,01000000,"&
"00000011,00000011,00000011,00000011,00000010,00000010,00000010,00000010,00000001,"&
"00000100,00000000,00000000,11110111,11111110,00000000,00000000,00000001,00000001,"&
"00000000,00000000,00000100,00000000,00000000,11100111,00000001,00000000,00000000,"&
"00000000,00000001,00000011,00000000,00000000,00000001,00000001,00000001,00000001,"&
"00000000,00000010,00000000,00000000,11111110,11111011,11111100,00000010,00000010,"&
"00000000,00000010,00000000,00000000,00000010,00000010,00000010,00000011,00000011,"&
"00000000,10110100,00000001,00000100,00000000,11111101,00000010,00000011,00000001,"&
"00000001,00000001,00000001,00000001,00000001,00000001,00000010,00000010,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000001,00000000,00000101,01000001,"&
"00000011,00000010,00000010,00000010,00000010,00000001,00000001,00000001,00000001,"&
"00000000,00000000,00000000,00000000,00000011,00000000,00000000,11000110,11110010,"&
"00000000,00000000,00000000,11000111,11110000,00000001,00000010,10100011,00000000,"&
"11111111,11000111,11101111,00000000,00000000,00000000,11111110,00001111,00000010,"&
"00000000,10100000,11111111,00000111,10011111,00000001,11110101,00000010,11111110,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"11111110,00000010,00000000,00000000,11111111,00000000,00000000,00000000,00000010,"&
"00000000,00000000,00000000,00000000,00000000,00000000,11111101,00000000,01000000,"&
"00000000,00000000,00000000,11111100,00000000,11111010,00000000,11111010,11100001,"&
"00011011,00000000,00000000,11100001,00000000,00000000,00000000,00000000,11111111,"&
"00000000,11100001,00000000,00010101,00000000,00000000,00110011,00001110,10110101,"&
"10111011,00000010,00000000,11111111,11110000,00110011,01000000,00000000,11000000,"&
"00000000,00000000,01000000,00000001,00000000,00000000,00000000,00000000,11111000,"&
"11001001,11001010,00000110,00000110,00000111,00000111,00000111,00000111,00000110,"&
"00000111,00000101,00000101,00000101,01000000,11010101,01000000,00000000,00000000,"&
"00000000,00000000,00000000,11001100,11010011,00000000,11001110,11010010,00000000,"&
"11010000,11010010,11010001,11010001,11010010,11010001,11010011,11010000,00000000,"&
"11010100,11001111,00000000,11010110,11001111,10110001,00000000,10110001,00000110,"&
"00010110,00001011,00000101,00011000,00000011,00000100,00100000,00000101,11110110,"&
"00100010,00000000,11011101,11001010,11110110,00000110,00100000,00000110,11110100,"&
"00000000,11011001,11001000,00000000,11000001,00000001,00000000,00000000,10110000,"&
"00000000,00000000,11100000,11000110,00000000,10111110,00000001,00000000,00000000,"&
"10101101,00000000,00000000,11001000,11101111,00000111,00001010,00000101,00000110,"&
"00100000,00000111,11101110,00000000,11011001,11000001,00000000,10111001,00000000,"&
"00000001,00000000,10101000,00000000,00000000,11100010,10111110,11101010,00000111,"&
"00001010,00000111,11101000,00000000,11011001,10111100,00000000,10110101,00000001,"&
"00000000,00000000,10100100,00000000,00000000,11100010,10111010,00000000,10110010,"&
"00000001,00000000,00000000,10100001,00000000,11100100,00000000,11010111,10110111,"&
"01000000,01000000,11100010,00000000,11011000,10110110,00110000,00110000,11100001,"&
"00000000,11011001,10110100,00000000,10101100,00000001,00000000,00000000,10011011,"&
"00000000,00000000,00000000,00000000,11011010,10110001,10010100,00000000,00000000,"&
"00000000,00000000,00000001,00001001,10010001,00000010,10010010,00111111,00000000,"&
"00000000,00000010,11100000,00000000,11111101,11111111,11111100,00000000,00001010,"&
"00000000,11011001,10101011,00000000,10100011,00000001,00000000,00000000,10010010,"&
"00000000,00000000,11011100,10101001,00000000,00000000,11010100,00000000,11011101,"&
"10100111,10001010,11111101,00000101,11010010,01000000,00000000,00111011,00111011,"&
"00000000,00000000,00000000,00000000,00000001,00000000,00000000,11000110,00001111,"&
"00000000,00000010,11010101,00000000,11111101,00000000,00000000,11011111,11100010,"&
"00000000,11011001,10100000,00000000,10011000,00000001,00000000,00000000,10000111,"&
"00000000,00000000,11100000,10011101,00000000,10010110,00000001,00000000,00000000,"&
"10000101,00000000,00000000,11100001,10011011,00000000,10010011,00000001,00000000,"&
"00000000,10000010,00001111,00000000,00000000,11111111,11000100,11111111,00000000,"&
"10110101,10111001,10111101,00111000,00000000,01111000,00000000,00000000,01001100,"&
"00000000,00110011,00110111,01100010,01100110,00000000,00100000,00110010,00000000,"&
"01010010,00100000,00100000,01110100,01100100,00101101,00001010,00000000,00101100,"&
"00100000,01100101,01010011,00101111,01110100,01000001,00000000,00101100,00100000,"&
"01101111,01100010,01110010,00000000,00101100,00100000,01110100,00000000,00100000,"&
"00100000,01100111,00100000,00100000,01010010,00000000,00100000,00100000,01100100,"&
"00000000,00100000,00100000,01101100,00000000,00100000,00100000,01100100,01110010,"&
"00000000,00100000,00100000,01110100,01101111,00000000,01001101,01101100,01100101,"&
"00000000,01000001,01100101,01110100,00000000,01100100,01110011,01100101,00000000,"&
"01101001,01100111,01110010,01101110,00100000,00110000,00111000,00101110,00000000,"&
"01101111,00000000,00100000,01100001,00000000,01101001,01110100,01000101,01001101,"&
"00000000,00100000,01100010,01110011,00000000,01101110,00100000,01111000,00000000,"&
"01110100,01101000,00111010,00000000,01111000,00000000,01110010,01101000,00111010,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,00000000,"&
"00000000,00000000,00000000,00000000,00000000,";




end package RAM_DATA;